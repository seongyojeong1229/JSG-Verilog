module xnor_gate_s(
    input a,
    input b,
    output y
    );

    xnor(y, a, b);

endmodule
