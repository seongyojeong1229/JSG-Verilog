module and_gate_s(
    input a,
    input b,
    output y
    );
    
    and(y,a,b);
    
endmodule
