module nor_gate_s(
    input a,
    input b,
    output y
    );

    nor(y, a, b);

endmodule
