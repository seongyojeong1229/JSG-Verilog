module xor_gate_s(
    input a,
    input b,
    output y
    );

    xor(y, a, b);

endmodule
