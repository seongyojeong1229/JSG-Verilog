module buffer_d(
    input a,
    output b
    );
    
    assign b = a;
    
endmodule
    
