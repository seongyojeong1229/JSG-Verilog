module buffer_s(
    input a,
    output b
    );
    
    buf(b,a);
    
endmodule
    
