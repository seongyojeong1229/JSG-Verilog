module not_gate_d(
    input a,
    output b
    );
    
    assign b = ~a;
endmodule

