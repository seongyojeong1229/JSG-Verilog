module not_gate_s(
    input a,
    output b
    );
    
    not(b,a);

endmodule

