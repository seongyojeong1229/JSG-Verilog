module nand_gate_s(
    input a,
    input b,
    output y
    );

    nand(y,a,b);

endmodule
