module or_gate_s(
    input a,
    input b,
    output y
    );

    or(y,a,b);
    
endmodule
